module();



endmodule
